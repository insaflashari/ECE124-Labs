 
LIBRARY ieee;
USE ieee.std_logic_1164.all; 
LIBRARY work;


ENTITY polarity_VHDL IS
	PORT (
			POLARITY_CONTRL, IN_1, IN_2, IN_3, IN_4: IN STD_LOGIC; 
			
			OUT_1, OUT_2, OUT_3, OUT_4: OUT STD_LOGIC
			);
			
END polarity_VHDL;

ARCHITECTURE simple_gates OF polarity_VHDL IS


BEGIN

OUT_1 <= POLARITY_CONTRL XNOR IN_1; 
OUT_2 <= POLARITY_CONTRL XNOR IN_2;
OUT_3 <= POLARITY_CONTRL XNOR IN_3;
OUT_4 <= POLARITY_CONTRL XNOR IN_4;

END simple_gates;